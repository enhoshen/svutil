// Copyright (C) Ganzin Technology - All Rights Reserved
// ---------------------------
// Unauthorized copying of this file, via any medium is strictly prohibited
// Proprietary and confidential
//
// Contributors
// ---------------------------
// En-Ho Shen <enhoshen@ganzin.com.tw>, 2020

`ifndef __DEFINE_SV__
`define __DEFINE_SV__

// packages

// sub-modules

`define D3 4

`endif //__DEFINE_SV__

