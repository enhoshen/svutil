`include "common/Define.sv"
`include "ValMatrix.sv"

