`include "Test.sv"

